magic
tech sky130A
timestamp 1743268417
<< nwell >>
rect -150 -50 1150 310
rect -150 -750 1150 -390
<< nmos >>
rect -35 -205 -20 -105
rect 315 -205 330 -105
rect 665 -205 680 -105
rect 1015 -205 1030 -105
rect -35 -905 -20 -805
rect 315 -905 330 -805
rect 665 -905 680 -805
rect 1015 -905 1030 -805
<< pmos >>
rect -35 -25 -20 175
rect 315 -25 330 175
rect 665 -25 680 175
rect 1015 -25 1030 175
rect -35 -725 -20 -525
rect 315 -725 330 -525
rect 665 -725 680 -525
rect 1015 -725 1030 -525
<< ndiff >>
rect -80 -115 -35 -105
rect -80 -135 -70 -115
rect -50 -135 -35 -115
rect -80 -175 -35 -135
rect -80 -195 -70 -175
rect -50 -195 -35 -175
rect -80 -205 -35 -195
rect -20 -115 25 -105
rect -20 -135 -5 -115
rect 15 -135 25 -115
rect -20 -175 25 -135
rect -20 -195 -5 -175
rect 15 -195 25 -175
rect -20 -205 25 -195
rect 270 -115 315 -105
rect 270 -135 280 -115
rect 300 -135 315 -115
rect 270 -175 315 -135
rect 270 -195 280 -175
rect 300 -195 315 -175
rect 270 -205 315 -195
rect 330 -115 375 -105
rect 330 -135 345 -115
rect 365 -135 375 -115
rect 330 -175 375 -135
rect 330 -195 345 -175
rect 365 -195 375 -175
rect 330 -205 375 -195
rect 620 -115 665 -105
rect 620 -135 630 -115
rect 650 -135 665 -115
rect 620 -175 665 -135
rect 620 -195 630 -175
rect 650 -195 665 -175
rect 620 -205 665 -195
rect 680 -115 725 -105
rect 680 -135 695 -115
rect 715 -135 725 -115
rect 680 -175 725 -135
rect 680 -195 695 -175
rect 715 -195 725 -175
rect 680 -205 725 -195
rect 970 -115 1015 -105
rect 970 -135 980 -115
rect 1000 -135 1015 -115
rect 970 -175 1015 -135
rect 970 -195 980 -175
rect 1000 -195 1015 -175
rect 970 -205 1015 -195
rect 1030 -115 1075 -105
rect 1030 -135 1045 -115
rect 1065 -135 1075 -115
rect 1030 -175 1075 -135
rect 1030 -195 1045 -175
rect 1065 -195 1075 -175
rect 1030 -205 1075 -195
rect -80 -815 -35 -805
rect -80 -835 -70 -815
rect -50 -835 -35 -815
rect -80 -875 -35 -835
rect -80 -895 -70 -875
rect -50 -895 -35 -875
rect -80 -905 -35 -895
rect -20 -815 25 -805
rect -20 -835 -5 -815
rect 15 -835 25 -815
rect -20 -875 25 -835
rect -20 -895 -5 -875
rect 15 -895 25 -875
rect -20 -905 25 -895
rect 270 -815 315 -805
rect 270 -835 280 -815
rect 300 -835 315 -815
rect 270 -875 315 -835
rect 270 -895 280 -875
rect 300 -895 315 -875
rect 270 -905 315 -895
rect 330 -815 375 -805
rect 330 -835 345 -815
rect 365 -835 375 -815
rect 330 -875 375 -835
rect 330 -895 345 -875
rect 365 -895 375 -875
rect 330 -905 375 -895
rect 620 -815 665 -805
rect 620 -835 630 -815
rect 650 -835 665 -815
rect 620 -875 665 -835
rect 620 -895 630 -875
rect 650 -895 665 -875
rect 620 -905 665 -895
rect 680 -815 725 -805
rect 680 -835 695 -815
rect 715 -835 725 -815
rect 680 -875 725 -835
rect 680 -895 695 -875
rect 715 -895 725 -875
rect 680 -905 725 -895
rect 970 -815 1015 -805
rect 970 -835 980 -815
rect 1000 -835 1015 -815
rect 970 -875 1015 -835
rect 970 -895 980 -875
rect 1000 -895 1015 -875
rect 970 -905 1015 -895
rect 1030 -815 1075 -805
rect 1030 -835 1045 -815
rect 1065 -835 1075 -815
rect 1030 -875 1075 -835
rect 1030 -895 1045 -875
rect 1065 -895 1075 -875
rect 1030 -905 1075 -895
<< pdiff >>
rect -80 165 -35 175
rect -80 145 -70 165
rect -50 145 -35 165
rect -80 90 -35 145
rect -80 70 -70 90
rect -50 70 -35 90
rect -80 5 -35 70
rect -80 -15 -70 5
rect -50 -15 -35 5
rect -80 -25 -35 -15
rect -20 165 25 175
rect -20 145 -5 165
rect 15 145 25 165
rect -20 90 25 145
rect -20 70 -5 90
rect 15 70 25 90
rect -20 5 25 70
rect -20 -15 -5 5
rect 15 -15 25 5
rect -20 -25 25 -15
rect 270 165 315 175
rect 270 145 280 165
rect 300 145 315 165
rect 270 90 315 145
rect 270 70 280 90
rect 300 70 315 90
rect 270 5 315 70
rect 270 -15 280 5
rect 300 -15 315 5
rect 270 -25 315 -15
rect 330 165 375 175
rect 330 145 345 165
rect 365 145 375 165
rect 330 90 375 145
rect 330 70 345 90
rect 365 70 375 90
rect 330 5 375 70
rect 330 -15 345 5
rect 365 -15 375 5
rect 330 -25 375 -15
rect 620 165 665 175
rect 620 145 630 165
rect 650 145 665 165
rect 620 90 665 145
rect 620 70 630 90
rect 650 70 665 90
rect 620 5 665 70
rect 620 -15 630 5
rect 650 -15 665 5
rect 620 -25 665 -15
rect 680 165 725 175
rect 680 145 695 165
rect 715 145 725 165
rect 680 90 725 145
rect 680 70 695 90
rect 715 70 725 90
rect 680 5 725 70
rect 680 -15 695 5
rect 715 -15 725 5
rect 680 -25 725 -15
rect 970 165 1015 175
rect 970 145 980 165
rect 1000 145 1015 165
rect 970 90 1015 145
rect 970 70 980 90
rect 1000 70 1015 90
rect 970 5 1015 70
rect 970 -15 980 5
rect 1000 -15 1015 5
rect 970 -25 1015 -15
rect 1030 165 1075 175
rect 1030 145 1045 165
rect 1065 145 1075 165
rect 1030 90 1075 145
rect 1030 70 1045 90
rect 1065 70 1075 90
rect 1030 5 1075 70
rect 1030 -15 1045 5
rect 1065 -15 1075 5
rect 1030 -25 1075 -15
rect -80 -535 -35 -525
rect -80 -555 -70 -535
rect -50 -555 -35 -535
rect -80 -610 -35 -555
rect -80 -630 -70 -610
rect -50 -630 -35 -610
rect -80 -695 -35 -630
rect -80 -715 -70 -695
rect -50 -715 -35 -695
rect -80 -725 -35 -715
rect -20 -535 25 -525
rect -20 -555 -5 -535
rect 15 -555 25 -535
rect -20 -610 25 -555
rect -20 -630 -5 -610
rect 15 -630 25 -610
rect -20 -695 25 -630
rect -20 -715 -5 -695
rect 15 -715 25 -695
rect -20 -725 25 -715
rect 270 -535 315 -525
rect 270 -555 280 -535
rect 300 -555 315 -535
rect 270 -610 315 -555
rect 270 -630 280 -610
rect 300 -630 315 -610
rect 270 -695 315 -630
rect 270 -715 280 -695
rect 300 -715 315 -695
rect 270 -725 315 -715
rect 330 -535 375 -525
rect 330 -555 345 -535
rect 365 -555 375 -535
rect 330 -610 375 -555
rect 330 -630 345 -610
rect 365 -630 375 -610
rect 330 -695 375 -630
rect 330 -715 345 -695
rect 365 -715 375 -695
rect 330 -725 375 -715
rect 620 -535 665 -525
rect 620 -555 630 -535
rect 650 -555 665 -535
rect 620 -610 665 -555
rect 620 -630 630 -610
rect 650 -630 665 -610
rect 620 -695 665 -630
rect 620 -715 630 -695
rect 650 -715 665 -695
rect 620 -725 665 -715
rect 680 -535 725 -525
rect 680 -555 695 -535
rect 715 -555 725 -535
rect 680 -610 725 -555
rect 680 -630 695 -610
rect 715 -630 725 -610
rect 680 -695 725 -630
rect 680 -715 695 -695
rect 715 -715 725 -695
rect 680 -725 725 -715
rect 970 -535 1015 -525
rect 970 -555 980 -535
rect 1000 -555 1015 -535
rect 970 -610 1015 -555
rect 970 -630 980 -610
rect 1000 -630 1015 -610
rect 970 -695 1015 -630
rect 970 -715 980 -695
rect 1000 -715 1015 -695
rect 970 -725 1015 -715
rect 1030 -535 1075 -525
rect 1030 -555 1045 -535
rect 1065 -555 1075 -535
rect 1030 -610 1075 -555
rect 1030 -630 1045 -610
rect 1065 -630 1075 -610
rect 1030 -695 1075 -630
rect 1030 -715 1045 -695
rect 1065 -715 1075 -695
rect 1030 -725 1075 -715
<< ndiffc >>
rect -70 -135 -50 -115
rect -70 -195 -50 -175
rect -5 -135 15 -115
rect -5 -195 15 -175
rect 280 -135 300 -115
rect 280 -195 300 -175
rect 345 -135 365 -115
rect 345 -195 365 -175
rect 630 -135 650 -115
rect 630 -195 650 -175
rect 695 -135 715 -115
rect 695 -195 715 -175
rect 980 -135 1000 -115
rect 980 -195 1000 -175
rect 1045 -135 1065 -115
rect 1045 -195 1065 -175
rect -70 -835 -50 -815
rect -70 -895 -50 -875
rect -5 -835 15 -815
rect -5 -895 15 -875
rect 280 -835 300 -815
rect 280 -895 300 -875
rect 345 -835 365 -815
rect 345 -895 365 -875
rect 630 -835 650 -815
rect 630 -895 650 -875
rect 695 -835 715 -815
rect 695 -895 715 -875
rect 980 -835 1000 -815
rect 980 -895 1000 -875
rect 1045 -835 1065 -815
rect 1045 -895 1065 -875
<< pdiffc >>
rect -70 145 -50 165
rect -70 70 -50 90
rect -70 -15 -50 5
rect -5 145 15 165
rect -5 70 15 90
rect -5 -15 15 5
rect 280 145 300 165
rect 280 70 300 90
rect 280 -15 300 5
rect 345 145 365 165
rect 345 70 365 90
rect 345 -15 365 5
rect 630 145 650 165
rect 630 70 650 90
rect 630 -15 650 5
rect 695 145 715 165
rect 695 70 715 90
rect 695 -15 715 5
rect 980 145 1000 165
rect 980 70 1000 90
rect 980 -15 1000 5
rect 1045 145 1065 165
rect 1045 70 1065 90
rect 1045 -15 1065 5
rect -70 -555 -50 -535
rect -70 -630 -50 -610
rect -70 -715 -50 -695
rect -5 -555 15 -535
rect -5 -630 15 -610
rect -5 -715 15 -695
rect 280 -555 300 -535
rect 280 -630 300 -610
rect 280 -715 300 -695
rect 345 -555 365 -535
rect 345 -630 365 -610
rect 345 -715 365 -695
rect 630 -555 650 -535
rect 630 -630 650 -610
rect 630 -715 650 -695
rect 695 -555 715 -535
rect 695 -630 715 -610
rect 695 -715 715 -695
rect 980 -555 1000 -535
rect 980 -630 1000 -610
rect 980 -715 1000 -695
rect 1045 -555 1065 -535
rect 1045 -630 1065 -610
rect 1045 -715 1065 -695
<< psubdiff >>
rect -80 -285 25 -270
rect -80 -305 -65 -285
rect -45 -305 -10 -285
rect 10 -305 25 -285
rect -80 -320 25 -305
rect 270 -285 375 -270
rect 270 -305 285 -285
rect 305 -305 340 -285
rect 360 -305 375 -285
rect 270 -320 375 -305
rect 620 -285 725 -270
rect 620 -305 635 -285
rect 655 -305 690 -285
rect 710 -305 725 -285
rect 620 -320 725 -305
rect 970 -285 1075 -270
rect 970 -305 985 -285
rect 1005 -305 1040 -285
rect 1060 -305 1075 -285
rect 970 -320 1075 -305
rect -80 -1015 25 -1000
rect -80 -1035 -65 -1015
rect -45 -1035 -10 -1015
rect 10 -1035 25 -1015
rect -80 -1050 25 -1035
rect 270 -1015 375 -1000
rect 270 -1035 285 -1015
rect 305 -1035 340 -1015
rect 360 -1035 375 -1015
rect 270 -1050 375 -1035
rect 620 -1015 725 -1000
rect 620 -1035 635 -1015
rect 655 -1035 690 -1015
rect 710 -1035 725 -1015
rect 620 -1050 725 -1035
rect 970 -1015 1075 -1000
rect 970 -1035 985 -1015
rect 1005 -1035 1040 -1015
rect 1060 -1035 1075 -1015
rect 970 -1050 1075 -1035
<< nsubdiff >>
rect -80 275 25 290
rect -80 255 -65 275
rect -45 255 -10 275
rect 10 255 25 275
rect -80 240 25 255
rect 270 275 375 290
rect 270 255 285 275
rect 305 255 340 275
rect 360 255 375 275
rect 270 240 375 255
rect 620 275 725 290
rect 620 255 635 275
rect 655 255 690 275
rect 710 255 725 275
rect 620 240 725 255
rect 970 275 1075 290
rect 970 255 985 275
rect 1005 255 1040 275
rect 1060 255 1075 275
rect 970 240 1075 255
rect -80 -425 25 -410
rect -80 -445 -65 -425
rect -45 -445 -10 -425
rect 10 -445 25 -425
rect -80 -460 25 -445
rect 270 -425 375 -410
rect 270 -445 285 -425
rect 305 -445 340 -425
rect 360 -445 375 -425
rect 270 -460 375 -445
rect 620 -425 725 -410
rect 620 -445 635 -425
rect 655 -445 690 -425
rect 710 -445 725 -425
rect 620 -460 725 -445
rect 970 -425 1075 -410
rect 970 -445 985 -425
rect 1005 -445 1040 -425
rect 1060 -445 1075 -425
rect 970 -460 1075 -445
<< psubdiffcont >>
rect -65 -305 -45 -285
rect -10 -305 10 -285
rect 285 -305 305 -285
rect 340 -305 360 -285
rect 635 -305 655 -285
rect 690 -305 710 -285
rect 985 -305 1005 -285
rect 1040 -305 1060 -285
rect -65 -1035 -45 -1015
rect -10 -1035 10 -1015
rect 285 -1035 305 -1015
rect 340 -1035 360 -1015
rect 635 -1035 655 -1015
rect 690 -1035 710 -1015
rect 985 -1035 1005 -1015
rect 1040 -1035 1060 -1015
<< nsubdiffcont >>
rect -65 255 -45 275
rect -10 255 10 275
rect 285 255 305 275
rect 340 255 360 275
rect 635 255 655 275
rect 690 255 710 275
rect 985 255 1005 275
rect 1040 255 1060 275
rect -65 -445 -45 -425
rect -10 -445 10 -425
rect 285 -445 305 -425
rect 340 -445 360 -425
rect 635 -445 655 -425
rect 690 -445 710 -425
rect 985 -445 1005 -425
rect 1040 -445 1060 -425
<< poly >>
rect 230 215 680 230
rect -35 175 -20 190
rect -35 -45 -20 -25
rect -70 -55 -20 -45
rect -70 -75 -60 -55
rect -40 -75 -20 -55
rect -70 -85 -20 -75
rect -35 -105 -20 -85
rect 165 -60 205 -50
rect 230 -60 245 215
rect 315 175 330 190
rect 665 175 680 215
rect 1015 175 1030 190
rect 315 -35 330 -25
rect 665 -35 680 -25
rect 1015 -35 1030 -25
rect 315 -50 505 -35
rect 665 -50 755 -35
rect 1015 -50 1145 -35
rect 165 -80 175 -60
rect 195 -80 245 -60
rect 490 -80 505 -50
rect 165 -90 205 -80
rect 230 -95 330 -80
rect 490 -95 680 -80
rect 315 -105 330 -95
rect 665 -105 680 -95
rect -35 -220 -20 -205
rect 315 -220 330 -205
rect 665 -230 680 -205
rect 455 -245 680 -230
rect 455 -315 470 -245
rect 445 -325 485 -315
rect 445 -345 455 -325
rect 475 -345 485 -325
rect 445 -355 485 -345
rect 35 -480 75 -470
rect 35 -485 45 -480
rect -35 -500 45 -485
rect 65 -500 75 -480
rect 455 -500 470 -355
rect 740 -500 755 -50
rect 1015 -105 1030 -90
rect 1015 -215 1030 -205
rect 1015 -230 1100 -215
rect 1085 -350 1100 -230
rect -35 -505 75 -500
rect -35 -525 -20 -505
rect 35 -510 75 -505
rect 315 -515 470 -500
rect 665 -515 755 -500
rect 840 -365 1100 -350
rect 1130 -355 1145 -50
rect 315 -525 330 -515
rect 665 -525 680 -515
rect -35 -745 -20 -725
rect -70 -755 -20 -745
rect 315 -735 330 -725
rect 665 -735 680 -725
rect 315 -750 505 -735
rect 665 -750 760 -735
rect -70 -775 -60 -755
rect -40 -775 -20 -755
rect -70 -785 -20 -775
rect -35 -805 -20 -785
rect 490 -780 505 -750
rect 315 -805 330 -790
rect 490 -795 680 -780
rect 665 -805 680 -795
rect -35 -920 -20 -905
rect 315 -945 330 -905
rect 665 -920 680 -905
rect 745 -945 760 -750
rect 315 -960 760 -945
rect 840 -965 855 -365
rect 1085 -500 1100 -365
rect 1125 -365 1165 -355
rect 1125 -385 1135 -365
rect 1155 -385 1165 -365
rect 1125 -395 1165 -385
rect 1015 -515 1100 -500
rect 1015 -525 1030 -515
rect 1015 -740 1030 -725
rect 1130 -780 1145 -395
rect 1015 -795 1145 -780
rect 1015 -805 1030 -795
rect 1015 -920 1030 -905
rect 835 -975 875 -965
rect 835 -995 845 -975
rect 865 -995 875 -975
rect 835 -1005 875 -995
<< polycont >>
rect -60 -75 -40 -55
rect 175 -80 195 -60
rect 455 -345 475 -325
rect 45 -500 65 -480
rect -60 -775 -40 -755
rect 1135 -385 1155 -365
rect 845 -995 865 -975
<< locali >>
rect -75 275 20 285
rect -75 255 -65 275
rect -45 255 -10 275
rect 10 255 20 275
rect -75 245 20 255
rect 275 275 370 285
rect 275 255 285 275
rect 305 255 340 275
rect 360 255 370 275
rect 275 245 370 255
rect 625 275 720 285
rect 625 255 635 275
rect 655 255 690 275
rect 710 255 720 275
rect 625 245 720 255
rect 975 275 1070 285
rect 975 255 985 275
rect 1005 255 1040 275
rect 1060 255 1070 275
rect 975 245 1070 255
rect -70 175 -50 245
rect 230 195 365 215
rect -80 165 -40 175
rect -80 145 -70 165
rect -50 145 -40 165
rect -80 90 -40 145
rect -80 70 -70 90
rect -50 70 -40 90
rect -80 5 -40 70
rect -80 -15 -70 5
rect -50 -15 -40 5
rect -80 -25 -40 -15
rect -15 165 25 175
rect -15 145 -5 165
rect 15 145 25 165
rect -15 90 25 145
rect -15 70 -5 90
rect 15 70 25 90
rect -15 5 25 70
rect -15 -15 -5 5
rect 15 -15 25 5
rect -15 -25 25 -15
rect -70 -55 -30 -45
rect -120 -75 -60 -55
rect -40 -75 -30 -55
rect -120 -335 -100 -75
rect -70 -85 -30 -75
rect -5 -60 15 -25
rect 165 -60 205 -50
rect -5 -80 175 -60
rect 195 -80 205 -60
rect -5 -105 15 -80
rect 165 -90 205 -80
rect -80 -115 -40 -105
rect -80 -135 -70 -115
rect -50 -135 -40 -115
rect -80 -175 -40 -135
rect -80 -195 -70 -175
rect -50 -195 -40 -175
rect -80 -205 -40 -195
rect -15 -115 25 -105
rect -15 -135 -5 -115
rect 15 -135 25 -115
rect 230 -115 250 195
rect 345 175 365 195
rect 580 195 715 215
rect 270 165 310 175
rect 270 145 280 165
rect 300 145 310 165
rect 270 90 310 145
rect 270 70 280 90
rect 300 70 310 90
rect 270 5 310 70
rect 270 -15 280 5
rect 300 -15 310 5
rect 270 -25 310 -15
rect 335 165 375 175
rect 335 145 345 165
rect 365 145 375 165
rect 335 90 375 145
rect 335 70 345 90
rect 365 70 375 90
rect 335 5 375 70
rect 335 -15 345 5
rect 365 -15 375 5
rect 335 -25 375 -15
rect 280 -50 300 -25
rect 280 -70 365 -50
rect 345 -105 365 -70
rect 270 -115 310 -105
rect 230 -135 280 -115
rect 300 -135 310 -115
rect -15 -175 25 -135
rect -15 -195 -5 -175
rect 15 -195 25 -175
rect -15 -205 25 -195
rect 270 -175 310 -135
rect 270 -195 280 -175
rect 300 -195 310 -175
rect 270 -205 310 -195
rect 335 -115 375 -105
rect 335 -135 345 -115
rect 365 -135 375 -115
rect 580 -115 600 195
rect 695 175 715 195
rect 930 195 1065 215
rect 620 165 660 175
rect 620 145 630 165
rect 650 145 660 165
rect 620 90 660 145
rect 620 70 630 90
rect 650 70 660 90
rect 620 5 660 70
rect 620 -15 630 5
rect 650 -15 660 5
rect 620 -25 660 -15
rect 685 165 725 175
rect 685 145 695 165
rect 715 145 725 165
rect 685 90 725 145
rect 685 70 695 90
rect 715 70 725 90
rect 685 5 725 70
rect 685 -15 695 5
rect 715 -15 725 5
rect 685 -25 725 -15
rect 630 -50 650 -25
rect 630 -70 715 -50
rect 695 -105 715 -70
rect 620 -115 660 -105
rect 580 -135 630 -115
rect 650 -135 660 -115
rect 335 -175 375 -135
rect 335 -195 345 -175
rect 365 -195 375 -175
rect 335 -205 375 -195
rect 620 -175 660 -135
rect 620 -195 630 -175
rect 650 -195 660 -175
rect 620 -205 660 -195
rect 685 -115 725 -105
rect 685 -135 695 -115
rect 715 -135 725 -115
rect 930 -115 950 195
rect 1045 175 1065 195
rect 970 165 1010 175
rect 970 145 980 165
rect 1000 145 1010 165
rect 970 90 1010 145
rect 970 70 980 90
rect 1000 70 1010 90
rect 970 5 1010 70
rect 970 -15 980 5
rect 1000 -15 1010 5
rect 970 -25 1010 -15
rect 1035 165 1075 175
rect 1035 145 1045 165
rect 1065 145 1075 165
rect 1035 90 1075 145
rect 1035 70 1045 90
rect 1065 70 1075 90
rect 1035 5 1075 70
rect 1035 -15 1045 5
rect 1065 -15 1075 5
rect 1035 -25 1075 -15
rect 980 -50 1000 -25
rect 980 -70 1065 -50
rect 1045 -105 1065 -70
rect 970 -115 1010 -105
rect 930 -135 980 -115
rect 1000 -135 1010 -115
rect 685 -175 725 -135
rect 685 -195 695 -175
rect 715 -195 725 -175
rect 685 -205 725 -195
rect 970 -175 1010 -135
rect 970 -195 980 -175
rect 1000 -195 1010 -175
rect 970 -205 1010 -195
rect 1035 -115 1075 -105
rect 1035 -135 1045 -115
rect 1065 -135 1075 -115
rect 1035 -175 1075 -135
rect 1035 -195 1045 -175
rect 1065 -195 1075 -175
rect 1035 -205 1075 -195
rect -70 -275 -50 -205
rect 280 -225 300 -205
rect 630 -225 650 -205
rect 1045 -225 1065 -205
rect 280 -245 1065 -225
rect -75 -285 20 -275
rect -75 -305 -65 -285
rect -45 -305 -10 -285
rect 10 -305 20 -285
rect -75 -315 20 -305
rect 275 -285 370 -275
rect 275 -305 285 -285
rect 305 -305 340 -285
rect 360 -305 370 -285
rect 275 -315 370 -305
rect 625 -285 720 -275
rect 625 -305 635 -285
rect 655 -305 690 -285
rect 710 -305 720 -285
rect 625 -315 720 -305
rect 975 -285 1070 -275
rect 975 -305 985 -285
rect 1005 -305 1040 -285
rect 1060 -305 1070 -285
rect 975 -315 1070 -305
rect 445 -325 485 -315
rect 445 -335 455 -325
rect -120 -345 455 -335
rect 475 -345 485 -325
rect -120 -355 485 -345
rect 1125 -365 1165 -355
rect 1125 -375 1135 -365
rect 110 -385 1135 -375
rect 1155 -385 1165 -365
rect 110 -395 1165 -385
rect -75 -425 20 -415
rect -75 -445 -65 -425
rect -45 -445 -10 -425
rect 10 -445 20 -425
rect -75 -455 20 -445
rect -70 -525 -50 -455
rect 35 -480 75 -470
rect 110 -480 130 -395
rect 275 -425 370 -415
rect 275 -445 285 -425
rect 305 -445 340 -425
rect 360 -445 370 -425
rect 275 -455 370 -445
rect 625 -425 720 -415
rect 625 -445 635 -425
rect 655 -445 690 -425
rect 710 -445 720 -425
rect 625 -455 720 -445
rect 975 -425 1070 -415
rect 975 -445 985 -425
rect 1005 -445 1040 -425
rect 1060 -445 1070 -425
rect 975 -455 1070 -445
rect 35 -500 45 -480
rect 65 -500 130 -480
rect 35 -510 75 -500
rect 230 -505 365 -485
rect -80 -535 -40 -525
rect -80 -555 -70 -535
rect -50 -555 -40 -535
rect -80 -610 -40 -555
rect -80 -630 -70 -610
rect -50 -630 -40 -610
rect -80 -695 -40 -630
rect -80 -715 -70 -695
rect -50 -715 -40 -695
rect -80 -725 -40 -715
rect -15 -535 25 -525
rect -15 -555 -5 -535
rect 15 -555 25 -535
rect -15 -610 25 -555
rect -15 -630 -5 -610
rect 15 -630 25 -610
rect -15 -695 25 -630
rect -15 -715 -5 -695
rect 15 -715 25 -695
rect -15 -725 25 -715
rect -70 -755 -30 -745
rect -70 -775 -60 -755
rect -40 -775 -30 -755
rect -70 -785 -30 -775
rect -5 -765 15 -725
rect -5 -785 85 -765
rect -5 -805 15 -785
rect -80 -815 -40 -805
rect -80 -835 -70 -815
rect -50 -835 -40 -815
rect -80 -875 -40 -835
rect -80 -895 -70 -875
rect -50 -895 -40 -875
rect -80 -905 -40 -895
rect -15 -815 25 -805
rect -15 -835 -5 -815
rect 15 -835 25 -815
rect -15 -875 25 -835
rect -15 -895 -5 -875
rect 15 -895 25 -875
rect -15 -905 25 -895
rect -70 -1005 -50 -905
rect 65 -965 85 -785
rect 230 -815 250 -505
rect 345 -525 365 -505
rect 580 -505 715 -485
rect 270 -535 310 -525
rect 270 -555 280 -535
rect 300 -555 310 -535
rect 270 -610 310 -555
rect 270 -630 280 -610
rect 300 -630 310 -610
rect 270 -695 310 -630
rect 270 -715 280 -695
rect 300 -715 310 -695
rect 270 -725 310 -715
rect 335 -535 375 -525
rect 335 -555 345 -535
rect 365 -555 375 -535
rect 335 -610 375 -555
rect 335 -630 345 -610
rect 365 -630 375 -610
rect 335 -695 375 -630
rect 335 -715 345 -695
rect 365 -715 375 -695
rect 335 -725 375 -715
rect 280 -755 300 -725
rect 280 -775 365 -755
rect 345 -805 365 -775
rect 270 -815 310 -805
rect 230 -835 280 -815
rect 300 -835 310 -815
rect 270 -875 310 -835
rect 270 -895 280 -875
rect 300 -895 310 -875
rect 270 -905 310 -895
rect 335 -815 375 -805
rect 335 -835 345 -815
rect 365 -835 375 -815
rect 580 -815 600 -505
rect 695 -525 715 -505
rect 930 -505 1065 -485
rect 620 -535 660 -525
rect 620 -555 630 -535
rect 650 -555 660 -535
rect 620 -610 660 -555
rect 620 -630 630 -610
rect 650 -630 660 -610
rect 620 -695 660 -630
rect 620 -715 630 -695
rect 650 -715 660 -695
rect 620 -725 660 -715
rect 685 -535 725 -525
rect 685 -555 695 -535
rect 715 -555 725 -535
rect 685 -610 725 -555
rect 685 -630 695 -610
rect 715 -630 725 -610
rect 685 -695 725 -630
rect 685 -715 695 -695
rect 715 -715 725 -695
rect 685 -725 725 -715
rect 630 -755 650 -725
rect 630 -775 715 -755
rect 695 -805 715 -775
rect 620 -815 660 -805
rect 580 -835 630 -815
rect 650 -835 660 -815
rect 335 -875 375 -835
rect 335 -895 345 -875
rect 365 -895 375 -875
rect 335 -905 375 -895
rect 620 -875 660 -835
rect 620 -895 630 -875
rect 650 -895 660 -875
rect 620 -905 660 -895
rect 685 -815 725 -805
rect 685 -835 695 -815
rect 715 -835 725 -815
rect 930 -815 950 -505
rect 1045 -525 1065 -505
rect 970 -535 1010 -525
rect 970 -555 980 -535
rect 1000 -555 1010 -535
rect 970 -610 1010 -555
rect 970 -630 980 -610
rect 1000 -630 1010 -610
rect 970 -695 1010 -630
rect 970 -715 980 -695
rect 1000 -715 1010 -695
rect 970 -725 1010 -715
rect 1035 -535 1075 -525
rect 1035 -555 1045 -535
rect 1065 -555 1075 -535
rect 1035 -610 1075 -555
rect 1035 -630 1045 -610
rect 1065 -630 1075 -610
rect 1035 -695 1075 -630
rect 1035 -715 1045 -695
rect 1065 -715 1075 -695
rect 1035 -725 1075 -715
rect 980 -755 1000 -725
rect 980 -775 1065 -755
rect 1045 -805 1065 -775
rect 970 -815 1010 -805
rect 930 -835 980 -815
rect 1000 -835 1010 -815
rect 685 -875 725 -835
rect 685 -895 695 -875
rect 715 -895 725 -875
rect 685 -905 725 -895
rect 970 -875 1010 -835
rect 970 -895 980 -875
rect 1000 -895 1010 -875
rect 970 -905 1010 -895
rect 1035 -815 1075 -805
rect 1035 -835 1045 -815
rect 1065 -835 1075 -815
rect 1035 -875 1075 -835
rect 1035 -895 1045 -875
rect 1065 -895 1075 -875
rect 1035 -905 1075 -895
rect 280 -925 300 -905
rect 630 -925 650 -905
rect 1045 -925 1065 -905
rect 280 -945 1065 -925
rect 65 -975 875 -965
rect 65 -985 845 -975
rect 835 -995 845 -985
rect 865 -995 875 -975
rect 835 -1005 875 -995
rect -75 -1015 20 -1005
rect -75 -1035 -65 -1015
rect -45 -1035 -10 -1015
rect 10 -1035 20 -1015
rect -75 -1045 20 -1035
rect 275 -1015 370 -1005
rect 275 -1035 285 -1015
rect 305 -1035 340 -1015
rect 360 -1035 370 -1015
rect 275 -1045 370 -1035
rect 625 -1015 720 -1005
rect 625 -1035 635 -1015
rect 655 -1035 690 -1015
rect 710 -1035 720 -1015
rect 625 -1045 720 -1035
rect 975 -1015 1070 -1005
rect 975 -1035 985 -1015
rect 1005 -1035 1040 -1015
rect 1060 -1035 1070 -1015
rect 975 -1045 1070 -1035
<< viali >>
rect -65 255 -45 275
rect -10 255 10 275
rect 285 255 305 275
rect 340 255 360 275
rect 635 255 655 275
rect 690 255 710 275
rect 985 255 1005 275
rect 1040 255 1060 275
rect -60 -75 -40 -55
rect 280 145 300 165
rect 630 70 650 90
rect 1045 -15 1065 5
rect -65 -305 -45 -285
rect -10 -305 10 -285
rect 285 -305 305 -285
rect 340 -305 360 -285
rect 635 -305 655 -285
rect 690 -305 710 -285
rect 985 -305 1005 -285
rect 1040 -305 1060 -285
rect -65 -445 -45 -425
rect -10 -445 10 -425
rect 285 -445 305 -425
rect 340 -445 360 -425
rect 635 -445 655 -425
rect 690 -445 710 -425
rect 985 -445 1005 -425
rect 1040 -445 1060 -425
rect -60 -775 -40 -755
rect 280 -555 300 -535
rect 630 -630 650 -610
rect 1045 -555 1065 -535
rect -65 -1035 -45 -1015
rect -10 -1035 10 -1015
rect 285 -1035 305 -1015
rect 340 -1035 360 -1015
rect 635 -1035 655 -1015
rect 690 -1035 710 -1015
rect 985 -1035 1005 -1015
rect 1040 -1035 1060 -1015
<< metal1 >>
rect -190 275 1190 285
rect -190 255 -65 275
rect -45 255 -10 275
rect 10 255 285 275
rect 305 255 340 275
rect 360 255 635 275
rect 655 255 690 275
rect 710 255 985 275
rect 1005 255 1040 275
rect 1060 255 1190 275
rect -190 245 1190 255
rect -190 165 310 175
rect -190 145 280 165
rect 300 145 310 165
rect -190 135 310 145
rect -190 90 660 100
rect -190 70 630 90
rect 650 70 660 90
rect -190 60 660 70
rect 1035 5 1245 15
rect 1035 -15 1045 5
rect 1065 -15 1245 5
rect 1035 -25 1245 -15
rect -190 -55 -30 -45
rect -190 -75 -60 -55
rect -40 -75 -30 -55
rect -190 -85 -30 -75
rect 1205 -275 1245 -25
rect -190 -285 1190 -275
rect -190 -305 -65 -285
rect -45 -305 -10 -285
rect 10 -305 285 -285
rect 305 -305 340 -285
rect 360 -305 635 -285
rect 655 -305 690 -285
rect 710 -305 985 -285
rect 1005 -305 1040 -285
rect 1060 -305 1190 -285
rect -190 -315 1190 -305
rect 1205 -315 1265 -275
rect -190 -425 1190 -415
rect -190 -445 -65 -425
rect -45 -445 -10 -425
rect 10 -445 285 -425
rect 305 -445 340 -425
rect 360 -445 635 -425
rect 655 -445 690 -425
rect 710 -445 985 -425
rect 1005 -445 1040 -425
rect 1060 -445 1190 -425
rect -190 -455 1190 -445
rect 1205 -525 1245 -315
rect -190 -535 310 -525
rect -190 -555 280 -535
rect 300 -555 310 -535
rect -190 -565 310 -555
rect 1035 -535 1245 -525
rect 1035 -555 1045 -535
rect 1065 -555 1245 -535
rect 1035 -565 1245 -555
rect -190 -610 660 -600
rect -190 -630 630 -610
rect 650 -630 660 -610
rect -190 -640 660 -630
rect -190 -755 -30 -745
rect -190 -775 -60 -755
rect -40 -775 -30 -755
rect -190 -785 -30 -775
rect -190 -1015 1190 -1005
rect -190 -1035 -65 -1015
rect -45 -1035 -10 -1015
rect 10 -1035 285 -1015
rect 305 -1035 340 -1015
rect 360 -1035 635 -1015
rect 655 -1035 690 -1015
rect 710 -1035 985 -1015
rect 1005 -1035 1040 -1015
rect 1060 -1035 1190 -1015
rect -190 -1045 1190 -1035
<< labels >>
rlabel metal1 -180 265 -180 265 1 vdd
rlabel metal1 -180 -435 -180 -435 1 vdd
rlabel metal1 -180 -295 -180 -295 1 gnd
rlabel metal1 1265 -315 1265 -275 7 output
rlabel metal1 -190 -85 -190 -45 3 s0
rlabel metal1 -190 -785 -190 -745 3 s1
rlabel metal1 -180 -1025 -180 -1025 1 gnd
rlabel metal1 -190 135 -190 175 3 I0
rlabel metal1 -190 60 -190 100 3 I1
rlabel metal1 -190 -565 -190 -525 3 I2
rlabel metal1 -190 -640 -190 -600 3 I3
<< end >>
